//`ifndef _DATAPATH_VH
//`define _DATAPATH_VH

localparam REG_IN_FROM_ACC = 1'b0;

localparam ACC_IN_FROM_IMM = 2'b00;
localparam ACC_IN_FROM_REG = 2'b01;
localparam ACC_IN_FROM_ALU = 2'b10;

//`endif
