localparam PC_FROM_REG   = 2'b00;
localparam PC_FROM_DATA  = 2'b01;
localparam PC_FROM_INST  = 2'b10;

